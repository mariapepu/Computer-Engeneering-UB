b = b+1/b